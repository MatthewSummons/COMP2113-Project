Save Exists
